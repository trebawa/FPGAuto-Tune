library verilog;
use verilog.vl_types.all;
entity nn_mult_test is
end nn_mult_test;
