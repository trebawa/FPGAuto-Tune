library verilog;
use verilog.vl_types.all;
entity main_fsm_test is
end main_fsm_test;
