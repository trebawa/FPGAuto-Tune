library verilog;
use verilog.vl_types.all;
entity serial_peak_finder is
    port(
        clk             : in     vl_logic;
        start           : in     vl_logic;
        data_in         : in     vl_logic_vector(31 downto 0);
        index           : in     vl_logic_vector(8 downto 0);
        peak_index      : out    vl_logic_vector(11 downto 0)
    );
end serial_peak_finder;
