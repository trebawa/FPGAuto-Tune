library verilog;
use verilog.vl_types.all;
entity peak_finder_test is
end peak_finder_test;
