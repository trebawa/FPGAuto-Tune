library verilog;
use verilog.vl_types.all;
entity note_lut is
    port(
        freq_fun        : in     vl_logic_vector(31 downto 0);
        note_name       : out    vl_logic_vector(3 downto 0);
        note_octave     : out    vl_logic_vector(2 downto 0);
        greater         : out    vl_logic
    );
end note_lut;
