library verilog;
use verilog.vl_types.all;
entity cordictest is
end cordictest;
