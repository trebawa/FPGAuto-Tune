library verilog;
use verilog.vl_types.all;
entity nn_multiplier_test is
end nn_multiplier_test;
