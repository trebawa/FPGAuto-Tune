library verilog;
use verilog.vl_types.all;
entity note_lut_test is
end note_lut_test;
