/*
    Automatic speech recognition processor (asrv2)

    Copyright 2014 MIT
    Author: Michael Price (pricem@mit.edu)
    
    Use and distribution of this code is restricted.
    See LICENSE file in top level project directory.
*/

/*
    Automatically generated code; please modify with care.
    File type: SROM
*/

module twiddle_lut #(
    parameter word_size = 36,
    parameter log_depth = 10,
    parameter use_compiled = 0
) (
    input clk,
    input reset,
    input [log_depth - 1 : 0] read_address,
    input read_enable,
    output reg read_valid,
    output reg [word_size - 1 : 0] read_data
);

generate if (use_compiled) begin: compiled_rom
    
    //	TODO: Add support for compiled ROM.
    
end
else begin: behav_rom
    reg [word_size - 1 : 0] out_reg;
    always @(*) read_data = out_reg;

    //	Synchronous assignment, real scalar
    always @(posedge clk) if (reset) begin
    	out_reg <= 0;
    end
    else begin
        read_valid <= read_enable;
    	if (read_enable) case (read_address)
    		//	36 bits
    		10'h000:	out_reg <= 36'h000010000; 
    		10'h001:	out_reg <= 36'hff9b8fffe; 
    		10'h002:	out_reg <= 36'hff370fffb; 
    		10'h003:	out_reg <= 36'hfed28fff4; 
    		10'h004:	out_reg <= 36'hfe6e0ffec; 
    		10'h005:	out_reg <= 36'hfe098ffe1; 
    		10'h006:	out_reg <= 36'hfda50ffd3; 
    		10'h007:	out_reg <= 36'hfd408ffc3; 
    		10'h008:	out_reg <= 36'hfcdc4ffb1; 
    		10'h009:	out_reg <= 36'hfc77cff9c; 
    		10'h00a:	out_reg <= 36'hfc138ff84; 
    		10'h00b:	out_reg <= 36'hfbaf0ff6a; 
    		10'h00c:	out_reg <= 36'hfb4acff4e; 
    		10'h00d:	out_reg <= 36'hfae68ff2f; 
    		10'h00e:	out_reg <= 36'hfa828ff0e; 
    		10'h00f:	out_reg <= 36'hfa1e4feea; 
    		10'h010:	out_reg <= 36'hf9ba4fec4; 
    		10'h011:	out_reg <= 36'hf9564fe9b; 
    		10'h012:	out_reg <= 36'hf8f24fe70; 
    		10'h013:	out_reg <= 36'hf88e4fe43; 
    		10'h014:	out_reg <= 36'hf82a8fe13; 
    		10'h015:	out_reg <= 36'hf7c6cfde0; 
    		10'h016:	out_reg <= 36'hf7634fdab; 
    		10'h017:	out_reg <= 36'hf6ff8fd74; 
    		10'h018:	out_reg <= 36'hf69c0fd3a; 
    		10'h019:	out_reg <= 36'hf638cfcfe; 
    		10'h01a:	out_reg <= 36'hf5d58fcbf; 
    		10'h01b:	out_reg <= 36'hf5724fc7e; 
    		10'h01c:	out_reg <= 36'hf50f0fc3b; 
    		10'h01d:	out_reg <= 36'hf4ac0fbf5; 
    		10'h01e:	out_reg <= 36'hf4494fbac; 
    		10'h01f:	out_reg <= 36'hf3e68fb61; 
    		10'h020:	out_reg <= 36'hf383cfb14; 
    		10'h021:	out_reg <= 36'hf3214fac5; 
    		10'h022:	out_reg <= 36'hf2becfa73; 
    		10'h023:	out_reg <= 36'hf25c8fa1e; 
    		10'h024:	out_reg <= 36'hf1fa4f9c7; 
    		10'h025:	out_reg <= 36'hf1984f96e; 
    		10'h026:	out_reg <= 36'hf1368f912; 
    		10'h027:	out_reg <= 36'hf0d4cf8b4; 
    		10'h028:	out_reg <= 36'hf0734f853; 
    		10'h029:	out_reg <= 36'hf011cf7f1; 
    		10'h02a:	out_reg <= 36'hefb08f78b; 
    		10'h02b:	out_reg <= 36'hef4f4f724; 
    		10'h02c:	out_reg <= 36'heeee4f6ba; 
    		10'h02d:	out_reg <= 36'hee8d8f64d; 
    		10'h02e:	out_reg <= 36'hee2ccf5de; 
    		10'h02f:	out_reg <= 36'hedcc8f56d; 
    		10'h030:	out_reg <= 36'hed6c0f4fa; 
    		10'h031:	out_reg <= 36'hed0c0f484; 
    		10'h032:	out_reg <= 36'hecac0f40b; 
    		10'h033:	out_reg <= 36'hec4c4f391; 
    		10'h034:	out_reg <= 36'hebeccf314; 
    		10'h035:	out_reg <= 36'heb8d8f294; 
    		10'h036:	out_reg <= 36'heb2e4f213; 
    		10'h037:	out_reg <= 36'heacf4f18f; 
    		10'h038:	out_reg <= 36'hea708f109; 
    		10'h039:	out_reg <= 36'hea120f080; 
    		10'h03a:	out_reg <= 36'he9b3ceff5; 
    		10'h03b:	out_reg <= 36'he9558ef68; 
    		10'h03c:	out_reg <= 36'he8f78eed8; 
    		10'h03d:	out_reg <= 36'he89a0ee46; 
    		10'h03e:	out_reg <= 36'he83c8edb2; 
    		10'h03f:	out_reg <= 36'he7df4ed1c; 
    		10'h040:	out_reg <= 36'he7824ec83; 
    		10'h041:	out_reg <= 36'he7258ebe8; 
    		10'h042:	out_reg <= 36'he6c90eb4b; 
    		10'h043:	out_reg <= 36'he66cceaab; 
    		10'h044:	out_reg <= 36'he610cea09; 
    		10'h045:	out_reg <= 36'he5b4ce965; 
    		10'h046:	out_reg <= 36'he5594e8bf; 
    		10'h047:	out_reg <= 36'he4fe0e816; 
    		10'h048:	out_reg <= 36'he4a30e76b; 
    		10'h049:	out_reg <= 36'he4484e6be; 
    		10'h04a:	out_reg <= 36'he3edce60f; 
    		10'h04b:	out_reg <= 36'he393ce55e; 
    		10'h04c:	out_reg <= 36'he339ce4aa; 
    		10'h04d:	out_reg <= 36'he2e00e3f4; 
    		10'h04e:	out_reg <= 36'he286ce33c; 
    		10'h04f:	out_reg <= 36'he22d8e282; 
    		10'h050:	out_reg <= 36'he1d4ce1c5; 
    		10'h051:	out_reg <= 36'he17c4e106; 
    		10'h052:	out_reg <= 36'he1240e046; 
    		10'h053:	out_reg <= 36'he0cc0df83; 
    		10'h054:	out_reg <= 36'he0748debe; 
    		10'h055:	out_reg <= 36'he01d4ddf6; 
    		10'h056:	out_reg <= 36'hdfc64dd2d; 
    		10'h057:	out_reg <= 36'hdf6f8dc61; 
    		10'h058:	out_reg <= 36'hdf190db94; 
    		10'h059:	out_reg <= 36'hdec30dac4; 
    		10'h05a:	out_reg <= 36'hde6d4d9f2; 
    		10'h05b:	out_reg <= 36'hde17cd91e; 
    		10'h05c:	out_reg <= 36'hddc2cd848; 
    		10'h05d:	out_reg <= 36'hdd6e0d770; 
    		10'h05e:	out_reg <= 36'hdd198d695; 
    		10'h05f:	out_reg <= 36'hdcc58d5b9; 
    		10'h060:	out_reg <= 36'hdc71cd4db; 
    		10'h061:	out_reg <= 36'hdc1e4d3fa; 
    		10'h062:	out_reg <= 36'hdbcb4d318; 
    		10'h063:	out_reg <= 36'hdb788d233; 
    		10'h064:	out_reg <= 36'hdb260d14d; 
    		10'h065:	out_reg <= 36'hdad40d064; 
    		10'h066:	out_reg <= 36'hda828cf7a; 
    		10'h067:	out_reg <= 36'hda310ce8d; 
    		10'h068:	out_reg <= 36'hd9e04cd9f; 
    		10'h069:	out_reg <= 36'hd98f8ccae; 
    		10'h06a:	out_reg <= 36'hd93f8cbbb; 
    		10'h06b:	out_reg <= 36'hd8ef8cac7; 
    		10'h06c:	out_reg <= 36'hd8a04c9d1; 
    		10'h06d:	out_reg <= 36'hd8510c8d8; 
    		10'h06e:	out_reg <= 36'hd8028c7de; 
    		10'h06f:	out_reg <= 36'hd7b44c6e2; 
    		10'h070:	out_reg <= 36'hd7664c5e4; 
    		10'h071:	out_reg <= 36'hd718cc4e3; 
    		10'h072:	out_reg <= 36'hd6cb8c3e2; 
    		10'h073:	out_reg <= 36'hd67ecc2de; 
    		10'h074:	out_reg <= 36'hd6328c1d8; 
    		10'h075:	out_reg <= 36'hd5e68c0d0; 
    		10'h076:	out_reg <= 36'hd59b0bfc7; 
    		10'h077:	out_reg <= 36'hd5500bebc; 
    		10'h078:	out_reg <= 36'hd5054bdae; 
    		10'h079:	out_reg <= 36'hd4bb0bca0; 
    		10'h07a:	out_reg <= 36'hd4714bb8f; 
    		10'h07b:	out_reg <= 36'hd427cba7c; 
    		10'h07c:	out_reg <= 36'hd3decb968; 
    		10'h07d:	out_reg <= 36'hd3960b852; 
    		10'h07e:	out_reg <= 36'hd34e0b73a; 
    		10'h07f:	out_reg <= 36'hd3064b620; 
    		10'h080:	out_reg <= 36'hd2bf0b504; 
    		10'h081:	out_reg <= 36'hd2780b3e7; 
    		10'h082:	out_reg <= 36'hd2318b2c8; 
    		10'h083:	out_reg <= 36'hd1eb8b1a8; 
    		10'h084:	out_reg <= 36'hd1a60b085; 
    		10'h085:	out_reg <= 36'hd1610af61; 
    		10'h086:	out_reg <= 36'hd11c4ae3b; 
    		10'h087:	out_reg <= 36'hd0d80ad14; 
    		10'h088:	out_reg <= 36'hd0948abeb; 
    		10'h089:	out_reg <= 36'hd0510aac0; 
    		10'h08a:	out_reg <= 36'hd00e4a994; 
    		10'h08b:	out_reg <= 36'hcfcc0a866; 
    		10'h08c:	out_reg <= 36'hcf8a0a736; 
    		10'h08d:	out_reg <= 36'hcf488a605; 
    		10'h08e:	out_reg <= 36'hcf078a4d2; 
    		10'h08f:	out_reg <= 36'hcec74a39d; 
    		10'h090:	out_reg <= 36'hce870a267; 
    		10'h091:	out_reg <= 36'hce478a12f; 
    		10'h092:	out_reg <= 36'hce0889ff6; 
    		10'h093:	out_reg <= 36'hcdca09ebc; 
    		10'h094:	out_reg <= 36'hcd8bc9d7f; 
    		10'h095:	out_reg <= 36'hcd4e49c42; 
    		10'h096:	out_reg <= 36'hcd1149b02; 
    		10'h097:	out_reg <= 36'hccd4899c2; 
    		10'h098:	out_reg <= 36'hcc984987f; 
    		10'h099:	out_reg <= 36'hcc5cc973c; 
    		10'h09a:	out_reg <= 36'hcc21895f6; 
    		10'h09b:	out_reg <= 36'hcbe7094b0; 
    		10'h09c:	out_reg <= 36'hcbacc9368; 
    		10'h09d:	out_reg <= 36'hcb734921e; 
    		10'h09e:	out_reg <= 36'hcb3a090d3; 
    		10'h09f:	out_reg <= 36'hcb0188f87; 
    		10'h0a0:	out_reg <= 36'hcac948e39; 
    		10'h0a1:	out_reg <= 36'hca91c8cea; 
    		10'h0a2:	out_reg <= 36'hca5ac8b9a; 
    		10'h0a3:	out_reg <= 36'hca2408a48; 
    		10'h0a4:	out_reg <= 36'hc9ee088f5; 
    		10'h0a5:	out_reg <= 36'hc9b8887a1; 
    		10'h0a6:	out_reg <= 36'hc9838864b; 
    		10'h0a7:	out_reg <= 36'hc94f084f4; 
    		10'h0a8:	out_reg <= 36'hc91b0839c; 
    		10'h0a9:	out_reg <= 36'hc8e7c8242; 
    		10'h0aa:	out_reg <= 36'hc8b4c80e7; 
    		10'h0ab:	out_reg <= 36'hc88287f8b; 
    		10'h0ac:	out_reg <= 36'hc85087e2e; 
    		10'h0ad:	out_reg <= 36'hc81f47cd0; 
    		10'h0ae:	out_reg <= 36'hc7ee87b70; 
    		10'h0af:	out_reg <= 36'hc7be87a0f; 
    		10'h0b0:	out_reg <= 36'hc78ec78ad; 
    		10'h0b1:	out_reg <= 36'hc75f8774a; 
    		10'h0b2:	out_reg <= 36'hc731075e5; 
    		10'h0b3:	out_reg <= 36'hc70307480; 
    		10'h0b4:	out_reg <= 36'hc6d587319; 
    		10'h0b5:	out_reg <= 36'hc6a8871b1; 
    		10'h0b6:	out_reg <= 36'hc67c47049; 
    		10'h0b7:	out_reg <= 36'hc65086edf; 
    		10'h0b8:	out_reg <= 36'hc62546d74; 
    		10'h0b9:	out_reg <= 36'hc5fa86c08; 
    		10'h0ba:	out_reg <= 36'hc5d046a9b; 
    		10'h0bb:	out_reg <= 36'hc5a6c692d; 
    		10'h0bc:	out_reg <= 36'hc57dc67bd; 
    		10'h0bd:	out_reg <= 36'hc5554664d; 
    		10'h0be:	out_reg <= 36'hc52d464dc; 
    		10'h0bf:	out_reg <= 36'hc5060636a; 
    		10'h0c0:	out_reg <= 36'hc4df461f7; 
    		10'h0c1:	out_reg <= 36'hc4b906083; 
    		10'h0c2:	out_reg <= 36'hc49385f0e; 
    		10'h0c3:	out_reg <= 36'hc46e85d98; 
    		10'h0c4:	out_reg <= 36'hc44a05c22; 
    		10'h0c5:	out_reg <= 36'hc42605aaa; 
    		10'h0c6:	out_reg <= 36'hc402c5931; 
    		10'h0c7:	out_reg <= 36'hc3e0057b8; 
    		10'h0c8:	out_reg <= 36'hc3bdc563e; 
    		10'h0c9:	out_reg <= 36'hc39c454c3; 
    		10'h0ca:	out_reg <= 36'hc37b45347; 
    		10'h0cb:	out_reg <= 36'hc35b051ca; 
    		10'h0cc:	out_reg <= 36'hc33b0504d; 
    		10'h0cd:	out_reg <= 36'hc31bc4ecf; 
    		10'h0ce:	out_reg <= 36'hc2fd44d50; 
    		10'h0cf:	out_reg <= 36'hc2df04bd0; 
    		10'h0d0:	out_reg <= 36'hc2c184a50; 
    		10'h0d1:	out_reg <= 36'hc2a4c48ce; 
    		10'h0d2:	out_reg <= 36'hc2888474d; 
    		10'h0d3:	out_reg <= 36'hc26cc45ca; 
    		10'h0d4:	out_reg <= 36'hc25184447; 
    		10'h0d5:	out_reg <= 36'hc237042c3; 
    		10'h0d6:	out_reg <= 36'hc21d4413e; 
    		10'h0d7:	out_reg <= 36'hc203c3fb9; 
    		10'h0d8:	out_reg <= 36'hc1eb43e33; 
    		10'h0d9:	out_reg <= 36'hc1d303cad; 
    		10'h0da:	out_reg <= 36'hc1bb83b26; 
    		10'h0db:	out_reg <= 36'hc1a48399f; 
    		10'h0dc:	out_reg <= 36'hc18e43817; 
    		10'h0dd:	out_reg <= 36'hc1788368e; 
    		10'h0de:	out_reg <= 36'hc16343505; 
    		10'h0df:	out_reg <= 36'hc14ec337b; 
    		10'h0e0:	out_reg <= 36'hc13b031f1; 
    		10'h0e1:	out_reg <= 36'hc127c3066; 
    		10'h0e2:	out_reg <= 36'hc11502edb; 
    		10'h0e3:	out_reg <= 36'hc102c2d50; 
    		10'h0e4:	out_reg <= 36'hc0f142bc4; 
    		10'h0e5:	out_reg <= 36'hc0e082a37; 
    		10'h0e6:	out_reg <= 36'hc0d0428aa; 
    		10'h0e7:	out_reg <= 36'hc0c08271d; 
    		10'h0e8:	out_reg <= 36'hc0b182590; 
    		10'h0e9:	out_reg <= 36'hc0a302402; 
    		10'h0ea:	out_reg <= 36'hc09542273; 
    		10'h0eb:	out_reg <= 36'hc088020e5; 
    		10'h0ec:	out_reg <= 36'hc07b41f56; 
    		10'h0ed:	out_reg <= 36'hc06f41dc7; 
    		10'h0ee:	out_reg <= 36'hc06401c37; 
    		10'h0ef:	out_reg <= 36'hc05941aa7; 
    		10'h0f0:	out_reg <= 36'hc04f01917; 
    		10'h0f1:	out_reg <= 36'hc04581787; 
    		10'h0f2:	out_reg <= 36'hc03c815f6; 
    		10'h0f3:	out_reg <= 36'hc03441466; 
    		10'h0f4:	out_reg <= 36'hc02c812d5; 
    		10'h0f5:	out_reg <= 36'hc02581144; 
    		10'h0f6:	out_reg <= 36'hc01f00fb2; 
    		10'h0f7:	out_reg <= 36'hc01900e21; 
    		10'h0f8:	out_reg <= 36'hc013c0c8f; 
    		10'h0f9:	out_reg <= 36'hc00f40afe; 
    		10'h0fa:	out_reg <= 36'hc00b4096c; 
    		10'h0fb:	out_reg <= 36'hc007c07da; 
    		10'h0fc:	out_reg <= 36'hc00500648; 
    		10'h0fd:	out_reg <= 36'hc003004b6; 
    		10'h0fe:	out_reg <= 36'hc00140324; 
    		10'h0ff:	out_reg <= 36'hc00080192; 
    		10'h100:	out_reg <= 36'hc00000000; 
    		10'h101:	out_reg <= 36'hc000bfe6e; 
    		10'h102:	out_reg <= 36'hc0017fcdc; 
    		10'h103:	out_reg <= 36'hc0033fb4a; 
    		10'h104:	out_reg <= 36'hc0053f9b8; 
    		10'h105:	out_reg <= 36'hc007ff826; 
    		10'h106:	out_reg <= 36'hc00b7f694; 
    		10'h107:	out_reg <= 36'hc00f7f502; 
    		10'h108:	out_reg <= 36'hc013ff371; 
    		10'h109:	out_reg <= 36'hc0193f1df; 
    		10'h10a:	out_reg <= 36'hc01f3f04e; 
    		10'h10b:	out_reg <= 36'hc025beebc; 
    		10'h10c:	out_reg <= 36'hc02cbed2b; 
    		10'h10d:	out_reg <= 36'hc0347eb9a; 
    		10'h10e:	out_reg <= 36'hc03cbea0a; 
    		10'h10f:	out_reg <= 36'hc045be879; 
    		10'h110:	out_reg <= 36'hc04f3e6e9; 
    		10'h111:	out_reg <= 36'hc0597e559; 
    		10'h112:	out_reg <= 36'hc0643e3c9; 
    		10'h113:	out_reg <= 36'hc06f7e239; 
    		10'h114:	out_reg <= 36'hc07b7e0aa; 
    		10'h115:	out_reg <= 36'hc0883df1b; 
    		10'h116:	out_reg <= 36'hc0957dd8d; 
    		10'h117:	out_reg <= 36'hc0a33dbfe; 
    		10'h118:	out_reg <= 36'hc0b1bda70; 
    		10'h119:	out_reg <= 36'hc0c0bd8e3; 
    		10'h11a:	out_reg <= 36'hc0d07d756; 
    		10'h11b:	out_reg <= 36'hc0e0bd5c9; 
    		10'h11c:	out_reg <= 36'hc0f17d43c; 
    		10'h11d:	out_reg <= 36'hc102fd2b0; 
    		10'h11e:	out_reg <= 36'hc1153d125; 
    		10'h11f:	out_reg <= 36'hc127fcf9a; 
    		10'h120:	out_reg <= 36'hc13b3ce0f; 
    		10'h121:	out_reg <= 36'hc14efcc85; 
    		10'h122:	out_reg <= 36'hc1637cafb; 
    		10'h123:	out_reg <= 36'hc178bc972; 
    		10'h124:	out_reg <= 36'hc18e7c7e9; 
    		10'h125:	out_reg <= 36'hc1a4bc661; 
    		10'h126:	out_reg <= 36'hc1bbbc4da; 
    		10'h127:	out_reg <= 36'hc1d33c353; 
    		10'h128:	out_reg <= 36'hc1eb7c1cd; 
    		10'h129:	out_reg <= 36'hc203fc047; 
    		10'h12a:	out_reg <= 36'hc21d7bec2; 
    		10'h12b:	out_reg <= 36'hc2373bd3d; 
    		10'h12c:	out_reg <= 36'hc251bbbb9; 
    		10'h12d:	out_reg <= 36'hc26cfba36; 
    		10'h12e:	out_reg <= 36'hc288bb8b3; 
    		10'h12f:	out_reg <= 36'hc2a4fb732; 
    		10'h130:	out_reg <= 36'hc2c1bb5b0; 
    		10'h131:	out_reg <= 36'hc2df3b430; 
    		10'h132:	out_reg <= 36'hc2fd7b2b0; 
    		10'h133:	out_reg <= 36'hc31bfb131; 
    		10'h134:	out_reg <= 36'hc33b3afb3; 
    		10'h135:	out_reg <= 36'hc35b3ae36; 
    		10'h136:	out_reg <= 36'hc37b7acb9; 
    		10'h137:	out_reg <= 36'hc39c7ab3d; 
    		10'h138:	out_reg <= 36'hc3bdfa9c2; 
    		10'h139:	out_reg <= 36'hc3e03a848; 
    		10'h13a:	out_reg <= 36'hc402fa6cf; 
    		10'h13b:	out_reg <= 36'hc4263a556; 
    		10'h13c:	out_reg <= 36'hc44a3a3de; 
    		10'h13d:	out_reg <= 36'hc46eba268; 
    		10'h13e:	out_reg <= 36'hc493ba0f2; 
    		10'h13f:	out_reg <= 36'hc4b939f7d; 
    		10'h140:	out_reg <= 36'hc4df79e09; 
    		10'h141:	out_reg <= 36'hc50639c96; 
    		10'h142:	out_reg <= 36'hc52d79b24; 
    		10'h143:	out_reg <= 36'hc555799b3; 
    		10'h144:	out_reg <= 36'hc57df9843; 
    		10'h145:	out_reg <= 36'hc5a6f96d3; 
    		10'h146:	out_reg <= 36'hc5d079565; 
    		10'h147:	out_reg <= 36'hc5fab93f8; 
    		10'h148:	out_reg <= 36'hc6257928c; 
    		10'h149:	out_reg <= 36'hc650b9121; 
    		10'h14a:	out_reg <= 36'hc67c78fb7; 
    		10'h14b:	out_reg <= 36'hc6a8b8e4f; 
    		10'h14c:	out_reg <= 36'hc6d5b8ce7; 
    		10'h14d:	out_reg <= 36'hc70338b80; 
    		10'h14e:	out_reg <= 36'hc73138a1b; 
    		10'h14f:	out_reg <= 36'hc75fb88b6; 
    		10'h150:	out_reg <= 36'hc78ef8753; 
    		10'h151:	out_reg <= 36'hc7beb85f1; 
    		10'h152:	out_reg <= 36'hc7eeb8490; 
    		10'h153:	out_reg <= 36'hc81f78330; 
    		10'h154:	out_reg <= 36'hc850b81d2; 
    		10'h155:	out_reg <= 36'hc882b8075; 
    		10'h156:	out_reg <= 36'hc8b4f7f19; 
    		10'h157:	out_reg <= 36'hc8e7f7dbe; 
    		10'h158:	out_reg <= 36'hc91b37c64; 
    		10'h159:	out_reg <= 36'hc94f37b0c; 
    		10'h15a:	out_reg <= 36'hc983b79b5; 
    		10'h15b:	out_reg <= 36'hc9b8b785f; 
    		10'h15c:	out_reg <= 36'hc9ee3770b; 
    		10'h15d:	out_reg <= 36'hca24375b8; 
    		10'h15e:	out_reg <= 36'hca5af7466; 
    		10'h15f:	out_reg <= 36'hca91f7316; 
    		10'h160:	out_reg <= 36'hcac9771c7; 
    		10'h161:	out_reg <= 36'hcb01b7079; 
    		10'h162:	out_reg <= 36'hcb3a36f2d; 
    		10'h163:	out_reg <= 36'hcb7376de2; 
    		10'h164:	out_reg <= 36'hcbacf6c98; 
    		10'h165:	out_reg <= 36'hcbe736b50; 
    		10'h166:	out_reg <= 36'hcc21b6a0a; 
    		10'h167:	out_reg <= 36'hcc5cf68c4; 
    		10'h168:	out_reg <= 36'hcc9876781; 
    		10'h169:	out_reg <= 36'hccd4b663e; 
    		10'h16a:	out_reg <= 36'hcd11764fe; 
    		10'h16b:	out_reg <= 36'hcd4e763be; 
    		10'h16c:	out_reg <= 36'hcd8bf6281; 
    		10'h16d:	out_reg <= 36'hcdca36144; 
    		10'h16e:	out_reg <= 36'hce08b600a; 
    		10'h16f:	out_reg <= 36'hce47b5ed1; 
    		10'h170:	out_reg <= 36'hce8735d99; 
    		10'h171:	out_reg <= 36'hcec775c63; 
    		10'h172:	out_reg <= 36'hcf07b5b2e; 
    		10'h173:	out_reg <= 36'hcf48b59fb; 
    		10'h174:	out_reg <= 36'hcf8a358ca; 
    		10'h175:	out_reg <= 36'hcfcc3579a; 
    		10'h176:	out_reg <= 36'hd00e7566c; 
    		10'h177:	out_reg <= 36'hd05135540; 
    		10'h178:	out_reg <= 36'hd094b5415; 
    		10'h179:	out_reg <= 36'hd0d8352ec; 
    		10'h17a:	out_reg <= 36'hd11c751c5; 
    		10'h17b:	out_reg <= 36'hd1613509f; 
    		10'h17c:	out_reg <= 36'hd1a634f7b; 
    		10'h17d:	out_reg <= 36'hd1ebb4e58; 
    		10'h17e:	out_reg <= 36'hd231b4d38; 
    		10'h17f:	out_reg <= 36'hd27834c19; 
    		10'h180:	out_reg <= 36'hd2bf34afc; 
    		10'h181:	out_reg <= 36'hd306749e0; 
    		10'h182:	out_reg <= 36'hd34e348c6; 
    		10'h183:	out_reg <= 36'hd396347ae; 
    		10'h184:	out_reg <= 36'hd3def4698; 
    		10'h185:	out_reg <= 36'hd427f4584; 
    		10'h186:	out_reg <= 36'hd47174471; 
    		10'h187:	out_reg <= 36'hd4bb34360; 
    		10'h188:	out_reg <= 36'hd50574252; 
    		10'h189:	out_reg <= 36'hd55034144; 
    		10'h18a:	out_reg <= 36'hd59b34039; 
    		10'h18b:	out_reg <= 36'hd5e6b3f30; 
    		10'h18c:	out_reg <= 36'hd632b3e28; 
    		10'h18d:	out_reg <= 36'hd67ef3d22; 
    		10'h18e:	out_reg <= 36'hd6cbb3c1e; 
    		10'h18f:	out_reg <= 36'hd718f3b1d; 
    		10'h190:	out_reg <= 36'hd76673a1c; 
    		10'h191:	out_reg <= 36'hd7b47391e; 
    		10'h192:	out_reg <= 36'hd802b3822; 
    		10'h193:	out_reg <= 36'hd85133728; 
    		10'h194:	out_reg <= 36'hd8a07362f; 
    		10'h195:	out_reg <= 36'hd8efb3539; 
    		10'h196:	out_reg <= 36'hd93fb3445; 
    		10'h197:	out_reg <= 36'hd98fb3352; 
    		10'h198:	out_reg <= 36'hd9e073261; 
    		10'h199:	out_reg <= 36'hda3133173; 
    		10'h19a:	out_reg <= 36'hda82b3086; 
    		10'h19b:	out_reg <= 36'hdad432f9c; 
    		10'h19c:	out_reg <= 36'hdb2632eb3; 
    		10'h19d:	out_reg <= 36'hdb78b2dcd; 
    		10'h19e:	out_reg <= 36'hdbcb72ce8; 
    		10'h19f:	out_reg <= 36'hdc1e72c06; 
    		10'h1a0:	out_reg <= 36'hdc71f2b25; 
    		10'h1a1:	out_reg <= 36'hdcc5b2a47; 
    		10'h1a2:	out_reg <= 36'hdd19b296b; 
    		10'h1a3:	out_reg <= 36'hdd6e32890; 
    		10'h1a4:	out_reg <= 36'hddc2f27b8; 
    		10'h1a5:	out_reg <= 36'hde17f26e2; 
    		10'h1a6:	out_reg <= 36'hde6d7260e; 
    		10'h1a7:	out_reg <= 36'hdec33253c; 
    		10'h1a8:	out_reg <= 36'hdf193246c; 
    		10'h1a9:	out_reg <= 36'hdf6fb239f; 
    		10'h1aa:	out_reg <= 36'hdfc6722d3; 
    		10'h1ab:	out_reg <= 36'he01d7220a; 
    		10'h1ac:	out_reg <= 36'he074b2142; 
    		10'h1ad:	out_reg <= 36'he0cc3207d; 
    		10'h1ae:	out_reg <= 36'he12431fba; 
    		10'h1af:	out_reg <= 36'he17c71efa; 
    		10'h1b0:	out_reg <= 36'he1d4f1e3b; 
    		10'h1b1:	out_reg <= 36'he22db1d7e; 
    		10'h1b2:	out_reg <= 36'he286f1cc4; 
    		10'h1b3:	out_reg <= 36'he2e031c0c; 
    		10'h1b4:	out_reg <= 36'he339f1b56; 
    		10'h1b5:	out_reg <= 36'he393f1aa2; 
    		10'h1b6:	out_reg <= 36'he3edf19f1; 
    		10'h1b7:	out_reg <= 36'he44871942; 
    		10'h1b8:	out_reg <= 36'he4a331895; 
    		10'h1b9:	out_reg <= 36'he4fe317ea; 
    		10'h1ba:	out_reg <= 36'he55971741; 
    		10'h1bb:	out_reg <= 36'he5b4f169b; 
    		10'h1bc:	out_reg <= 36'he610f15f7; 
    		10'h1bd:	out_reg <= 36'he66cf1555; 
    		10'h1be:	out_reg <= 36'he6c9314b5; 
    		10'h1bf:	out_reg <= 36'he725b1418; 
    		10'h1c0:	out_reg <= 36'he7827137d; 
    		10'h1c1:	out_reg <= 36'he7df712e4; 
    		10'h1c2:	out_reg <= 36'he83cb124e; 
    		10'h1c3:	out_reg <= 36'he89a311ba; 
    		10'h1c4:	out_reg <= 36'he8f7b1128; 
    		10'h1c5:	out_reg <= 36'he955b1098; 
    		10'h1c6:	out_reg <= 36'he9b3f100b; 
    		10'h1c7:	out_reg <= 36'hea1230f80; 
    		10'h1c8:	out_reg <= 36'hea70b0ef7; 
    		10'h1c9:	out_reg <= 36'heacf70e71; 
    		10'h1ca:	out_reg <= 36'heb2e70ded; 
    		10'h1cb:	out_reg <= 36'heb8db0d6c; 
    		10'h1cc:	out_reg <= 36'hebecf0cec; 
    		10'h1cd:	out_reg <= 36'hec4c70c6f; 
    		10'h1ce:	out_reg <= 36'hecac30bf5; 
    		10'h1cf:	out_reg <= 36'hed0c30b7c; 
    		10'h1d0:	out_reg <= 36'hed6c30b06; 
    		10'h1d1:	out_reg <= 36'hedccb0a93; 
    		10'h1d2:	out_reg <= 36'hee2cf0a22; 
    		10'h1d3:	out_reg <= 36'hee8db09b3; 
    		10'h1d4:	out_reg <= 36'heeee70946; 
    		10'h1d5:	out_reg <= 36'hef4f708dc; 
    		10'h1d6:	out_reg <= 36'hefb0b0875; 
    		10'h1d7:	out_reg <= 36'hf011f080f; 
    		10'h1d8:	out_reg <= 36'hf073707ad; 
    		10'h1d9:	out_reg <= 36'hf0d4f074c; 
    		10'h1da:	out_reg <= 36'hf136b06ee; 
    		10'h1db:	out_reg <= 36'hf19870692; 
    		10'h1dc:	out_reg <= 36'hf1fa70639; 
    		10'h1dd:	out_reg <= 36'hf25cb05e2; 
    		10'h1de:	out_reg <= 36'hf2bef058d; 
    		10'h1df:	out_reg <= 36'hf3217053b; 
    		10'h1e0:	out_reg <= 36'hf383f04ec; 
    		10'h1e1:	out_reg <= 36'hf3e6b049f; 
    		10'h1e2:	out_reg <= 36'hf44970454; 
    		10'h1e3:	out_reg <= 36'hf4ac3040b; 
    		10'h1e4:	out_reg <= 36'hf50f303c5; 
    		10'h1e5:	out_reg <= 36'hf57270382; 
    		10'h1e6:	out_reg <= 36'hf5d5b0341; 
    		10'h1e7:	out_reg <= 36'hf638f0302; 
    		10'h1e8:	out_reg <= 36'hf69c302c6; 
    		10'h1e9:	out_reg <= 36'hf6ffb028c; 
    		10'h1ea:	out_reg <= 36'hf76370255; 
    		10'h1eb:	out_reg <= 36'hf7c6f0220; 
    		10'h1ec:	out_reg <= 36'hf82ab01ed; 
    		10'h1ed:	out_reg <= 36'hf88e701bd; 
    		10'h1ee:	out_reg <= 36'hf8f270190; 
    		10'h1ef:	out_reg <= 36'hf95670165; 
    		10'h1f0:	out_reg <= 36'hf9ba7013c; 
    		10'h1f1:	out_reg <= 36'hfa1e70116; 
    		10'h1f2:	out_reg <= 36'hfa82b00f2; 
    		10'h1f3:	out_reg <= 36'hfae6b00d1; 
    		10'h1f4:	out_reg <= 36'hfb4af00b2; 
    		10'h1f5:	out_reg <= 36'hfbaf30096; 
    		10'h1f6:	out_reg <= 36'hfc13b007c; 
    		10'h1f7:	out_reg <= 36'hfc77f0064; 
    		10'h1f8:	out_reg <= 36'hfcdc7004f; 
    		10'h1f9:	out_reg <= 36'hfd40b003d; 
    		10'h1fa:	out_reg <= 36'hfda53002d; 
    		10'h1fb:	out_reg <= 36'hfe09b001f; 
    		10'h1fc:	out_reg <= 36'hfe6e30014; 
    		10'h1fd:	out_reg <= 36'hfed2b000c; 
    		10'h1fe:	out_reg <= 36'hff3730005; 
    		10'h1ff:	out_reg <= 36'hff9bb0002; 
    		10'h200:	out_reg <= 36'h000030000; 
    		10'h201:	out_reg <= 36'h0064b0002; 
    		10'h202:	out_reg <= 36'h00c930005; 
    		10'h203:	out_reg <= 36'h012db000c; 
    		10'h204:	out_reg <= 36'h019230014; 
    		10'h205:	out_reg <= 36'h01f6b001f; 
    		10'h206:	out_reg <= 36'h025b3002d; 
    		10'h207:	out_reg <= 36'h02bfb003d; 
    		10'h208:	out_reg <= 36'h0323f004f; 
    		10'h209:	out_reg <= 36'h038870064; 
    		10'h20a:	out_reg <= 36'h03ecb007c; 
    		10'h20b:	out_reg <= 36'h045130096; 
    		10'h20c:	out_reg <= 36'h04b5700b2; 
    		10'h20d:	out_reg <= 36'h0519b00d1; 
    		10'h20e:	out_reg <= 36'h057db00f2; 
    		10'h20f:	out_reg <= 36'h05e1f0116; 
    		10'h210:	out_reg <= 36'h0645f013c; 
    		10'h211:	out_reg <= 36'h06a9f0165; 
    		10'h212:	out_reg <= 36'h070df0190; 
    		10'h213:	out_reg <= 36'h0771f01bd; 
    		10'h214:	out_reg <= 36'h07d5b01ed; 
    		10'h215:	out_reg <= 36'h083970220; 
    		10'h216:	out_reg <= 36'h089cf0255; 
    		10'h217:	out_reg <= 36'h0900b028c; 
    		10'h218:	out_reg <= 36'h0964302c6; 
    		10'h219:	out_reg <= 36'h09c770302; 
    		10'h21a:	out_reg <= 36'h0a2ab0341; 
    		10'h21b:	out_reg <= 36'h0a8df0382; 
    		10'h21c:	out_reg <= 36'h0af1303c5; 
    		10'h21d:	out_reg <= 36'h0b543040b; 
    		10'h21e:	out_reg <= 36'h0bb6f0454; 
    		10'h21f:	out_reg <= 36'h0c19b049f; 
    		10'h220:	out_reg <= 36'h0c7c704ec; 
    		10'h221:	out_reg <= 36'h0cdef053b; 
    		10'h222:	out_reg <= 36'h0d417058d; 
    		10'h223:	out_reg <= 36'h0da3b05e2; 
    		10'h224:	out_reg <= 36'h0e05f0639; 
    		10'h225:	out_reg <= 36'h0e67f0692; 
    		10'h226:	out_reg <= 36'h0ec9b06ee; 
    		10'h227:	out_reg <= 36'h0f2b7074c; 
    		10'h228:	out_reg <= 36'h0f8cf07ad; 
    		10'h229:	out_reg <= 36'h0fee7080f; 
    		10'h22a:	out_reg <= 36'h104fb0875; 
    		10'h22b:	out_reg <= 36'h10b0f08dc; 
    		10'h22c:	out_reg <= 36'h1111f0946; 
    		10'h22d:	out_reg <= 36'h1172b09b3; 
    		10'h22e:	out_reg <= 36'h11d370a22; 
    		10'h22f:	out_reg <= 36'h1233b0a93; 
    		10'h230:	out_reg <= 36'h129430b06; 
    		10'h231:	out_reg <= 36'h12f430b7c; 
    		10'h232:	out_reg <= 36'h135430bf5; 
    		10'h233:	out_reg <= 36'h13b3f0c6f; 
    		10'h234:	out_reg <= 36'h141370cec; 
    		10'h235:	out_reg <= 36'h1472b0d6c; 
    		10'h236:	out_reg <= 36'h14d1f0ded; 
    		10'h237:	out_reg <= 36'h1530f0e71; 
    		10'h238:	out_reg <= 36'h158fb0ef7; 
    		10'h239:	out_reg <= 36'h15ee30f80; 
    		10'h23a:	out_reg <= 36'h164c7100b; 
    		10'h23b:	out_reg <= 36'h16aab1098; 
    		10'h23c:	out_reg <= 36'h1708b1128; 
    		10'h23d:	out_reg <= 36'h1766311ba; 
    		10'h23e:	out_reg <= 36'h17c3b124e; 
    		10'h23f:	out_reg <= 36'h1820f12e4; 
    		10'h240:	out_reg <= 36'h187df137d; 
    		10'h241:	out_reg <= 36'h18dab1418; 
    		10'h242:	out_reg <= 36'h1937314b5; 
    		10'h243:	out_reg <= 36'h199371555; 
    		10'h244:	out_reg <= 36'h19ef715f7; 
    		10'h245:	out_reg <= 36'h1a4b7169b; 
    		10'h246:	out_reg <= 36'h1aa6f1741; 
    		10'h247:	out_reg <= 36'h1b02317ea; 
    		10'h248:	out_reg <= 36'h1b5d31895; 
    		10'h249:	out_reg <= 36'h1bb7f1942; 
    		10'h24a:	out_reg <= 36'h1c12719f1; 
    		10'h24b:	out_reg <= 36'h1c6c71aa2; 
    		10'h24c:	out_reg <= 36'h1cc671b56; 
    		10'h24d:	out_reg <= 36'h1d2031c0c; 
    		10'h24e:	out_reg <= 36'h1d7971cc4; 
    		10'h24f:	out_reg <= 36'h1dd2b1d7e; 
    		10'h250:	out_reg <= 36'h1e2b71e3b; 
    		10'h251:	out_reg <= 36'h1e83f1efa; 
    		10'h252:	out_reg <= 36'h1edc31fba; 
    		10'h253:	out_reg <= 36'h1f343207d; 
    		10'h254:	out_reg <= 36'h1f8bb2142; 
    		10'h255:	out_reg <= 36'h1fe2f220a; 
    		10'h256:	out_reg <= 36'h2039f22d3; 
    		10'h257:	out_reg <= 36'h2090b239f; 
    		10'h258:	out_reg <= 36'h20e73246c; 
    		10'h259:	out_reg <= 36'h213d3253c; 
    		10'h25a:	out_reg <= 36'h2192f260e; 
    		10'h25b:	out_reg <= 36'h21e8726e2; 
    		10'h25c:	out_reg <= 36'h223d727b8; 
    		10'h25d:	out_reg <= 36'h229232890; 
    		10'h25e:	out_reg <= 36'h22e6b296b; 
    		10'h25f:	out_reg <= 36'h233ab2a47; 
    		10'h260:	out_reg <= 36'h238e72b25; 
    		10'h261:	out_reg <= 36'h23e1f2c06; 
    		10'h262:	out_reg <= 36'h2434f2ce8; 
    		10'h263:	out_reg <= 36'h2487b2dcd; 
    		10'h264:	out_reg <= 36'h24da32eb3; 
    		10'h265:	out_reg <= 36'h252c32f9c; 
    		10'h266:	out_reg <= 36'h257db3086; 
    		10'h267:	out_reg <= 36'h25cf33173; 
    		10'h268:	out_reg <= 36'h261ff3261; 
    		10'h269:	out_reg <= 36'h2670b3352; 
    		10'h26a:	out_reg <= 36'h26c0b3445; 
    		10'h26b:	out_reg <= 36'h2710b3539; 
    		10'h26c:	out_reg <= 36'h275ff362f; 
    		10'h26d:	out_reg <= 36'h27af33728; 
    		10'h26e:	out_reg <= 36'h27fdb3822; 
    		10'h26f:	out_reg <= 36'h284bf391e; 
    		10'h270:	out_reg <= 36'h2899f3a1c; 
    		10'h271:	out_reg <= 36'h28e773b1d; 
    		10'h272:	out_reg <= 36'h2934b3c1e; 
    		10'h273:	out_reg <= 36'h298173d22; 
    		10'h274:	out_reg <= 36'h29cdb3e28; 
    		10'h275:	out_reg <= 36'h2a19b3f30; 
    		10'h276:	out_reg <= 36'h2a6534039; 
    		10'h277:	out_reg <= 36'h2ab034144; 
    		10'h278:	out_reg <= 36'h2afaf4252; 
    		10'h279:	out_reg <= 36'h2b4534360; 
    		10'h27a:	out_reg <= 36'h2b8ef4471; 
    		10'h27b:	out_reg <= 36'h2bd874584; 
    		10'h27c:	out_reg <= 36'h2c2174698; 
    		10'h27d:	out_reg <= 36'h2c6a347ae; 
    		10'h27e:	out_reg <= 36'h2cb2348c6; 
    		10'h27f:	out_reg <= 36'h2cf9f49e0; 
    		10'h280:	out_reg <= 36'h2d4134afc; 
    		10'h281:	out_reg <= 36'h2d8834c19; 
    		10'h282:	out_reg <= 36'h2dceb4d38; 
    		10'h283:	out_reg <= 36'h2e14b4e58; 
    		10'h284:	out_reg <= 36'h2e5a34f7b; 
    		10'h285:	out_reg <= 36'h2e9f3509f; 
    		10'h286:	out_reg <= 36'h2ee3f51c5; 
    		10'h287:	out_reg <= 36'h2f28352ec; 
    		10'h288:	out_reg <= 36'h2f6bb5415; 
    		10'h289:	out_reg <= 36'h2faf35540; 
    		10'h28a:	out_reg <= 36'h2ff1f566c; 
    		10'h28b:	out_reg <= 36'h30343579a; 
    		10'h28c:	out_reg <= 36'h3076358ca; 
    		10'h28d:	out_reg <= 36'h30b7b59fb; 
    		10'h28e:	out_reg <= 36'h30f8b5b2e; 
    		10'h28f:	out_reg <= 36'h3138f5c63; 
    		10'h290:	out_reg <= 36'h317935d99; 
    		10'h291:	out_reg <= 36'h31b8b5ed1; 
    		10'h292:	out_reg <= 36'h31f7b600a; 
    		10'h293:	out_reg <= 36'h323636144; 
    		10'h294:	out_reg <= 36'h327476281; 
    		10'h295:	out_reg <= 36'h32b1f63be; 
    		10'h296:	out_reg <= 36'h32eef64fe; 
    		10'h297:	out_reg <= 36'h332bb663e; 
    		10'h298:	out_reg <= 36'h3367f6781; 
    		10'h299:	out_reg <= 36'h33a3768c4; 
    		10'h29a:	out_reg <= 36'h33deb6a0a; 
    		10'h29b:	out_reg <= 36'h341936b50; 
    		10'h29c:	out_reg <= 36'h345376c98; 
    		10'h29d:	out_reg <= 36'h348cf6de2; 
    		10'h29e:	out_reg <= 36'h34c636f2d; 
    		10'h29f:	out_reg <= 36'h34feb7079; 
    		10'h2a0:	out_reg <= 36'h3536f71c7; 
    		10'h2a1:	out_reg <= 36'h356e77316; 
    		10'h2a2:	out_reg <= 36'h35a577466; 
    		10'h2a3:	out_reg <= 36'h35dc375b8; 
    		10'h2a4:	out_reg <= 36'h36123770b; 
    		10'h2a5:	out_reg <= 36'h3647b785f; 
    		10'h2a6:	out_reg <= 36'h367cb79b5; 
    		10'h2a7:	out_reg <= 36'h36b137b0c; 
    		10'h2a8:	out_reg <= 36'h36e537c64; 
    		10'h2a9:	out_reg <= 36'h371877dbe; 
    		10'h2aa:	out_reg <= 36'h374b77f19; 
    		10'h2ab:	out_reg <= 36'h377db8075; 
    		10'h2ac:	out_reg <= 36'h37afb81d2; 
    		10'h2ad:	out_reg <= 36'h37e0f8330; 
    		10'h2ae:	out_reg <= 36'h3811b8490; 
    		10'h2af:	out_reg <= 36'h3841b85f1; 
    		10'h2b0:	out_reg <= 36'h387178753; 
    		10'h2b1:	out_reg <= 36'h38a0b88b6; 
    		10'h2b2:	out_reg <= 36'h38cf38a1b; 
    		10'h2b3:	out_reg <= 36'h38fd38b80; 
    		10'h2b4:	out_reg <= 36'h392ab8ce7; 
    		10'h2b5:	out_reg <= 36'h3957b8e4f; 
    		10'h2b6:	out_reg <= 36'h3983f8fb7; 
    		10'h2b7:	out_reg <= 36'h39afb9121; 
    		10'h2b8:	out_reg <= 36'h39daf928c; 
    		10'h2b9:	out_reg <= 36'h3a05b93f8; 
    		10'h2ba:	out_reg <= 36'h3a2ff9565; 
    		10'h2bb:	out_reg <= 36'h3a59796d3; 
    		10'h2bc:	out_reg <= 36'h3a8279843; 
    		10'h2bd:	out_reg <= 36'h3aaaf99b3; 
    		10'h2be:	out_reg <= 36'h3ad2f9b24; 
    		10'h2bf:	out_reg <= 36'h3afa39c96; 
    		10'h2c0:	out_reg <= 36'h3b20f9e09; 
    		10'h2c1:	out_reg <= 36'h3b4739f7d; 
    		10'h2c2:	out_reg <= 36'h3b6cba0f2; 
    		10'h2c3:	out_reg <= 36'h3b91ba268; 
    		10'h2c4:	out_reg <= 36'h3bb63a3de; 
    		10'h2c5:	out_reg <= 36'h3bda3a556; 
    		10'h2c6:	out_reg <= 36'h3bfd7a6cf; 
    		10'h2c7:	out_reg <= 36'h3c203a848; 
    		10'h2c8:	out_reg <= 36'h3c427a9c2; 
    		10'h2c9:	out_reg <= 36'h3c63fab3d; 
    		10'h2ca:	out_reg <= 36'h3c84facb9; 
    		10'h2cb:	out_reg <= 36'h3ca53ae36; 
    		10'h2cc:	out_reg <= 36'h3cc53afb3; 
    		10'h2cd:	out_reg <= 36'h3ce47b131; 
    		10'h2ce:	out_reg <= 36'h3d02fb2b0; 
    		10'h2cf:	out_reg <= 36'h3d213b430; 
    		10'h2d0:	out_reg <= 36'h3d3ebb5b0; 
    		10'h2d1:	out_reg <= 36'h3d5b7b732; 
    		10'h2d2:	out_reg <= 36'h3d77bb8b3; 
    		10'h2d3:	out_reg <= 36'h3d937ba36; 
    		10'h2d4:	out_reg <= 36'h3daebbbb9; 
    		10'h2d5:	out_reg <= 36'h3dc93bd3d; 
    		10'h2d6:	out_reg <= 36'h3de2fbec2; 
    		10'h2d7:	out_reg <= 36'h3dfc7c047; 
    		10'h2d8:	out_reg <= 36'h3e14fc1cd; 
    		10'h2d9:	out_reg <= 36'h3e2d3c353; 
    		10'h2da:	out_reg <= 36'h3e44bc4da; 
    		10'h2db:	out_reg <= 36'h3e5bbc661; 
    		10'h2dc:	out_reg <= 36'h3e71fc7e9; 
    		10'h2dd:	out_reg <= 36'h3e87bc972; 
    		10'h2de:	out_reg <= 36'h3e9cfcafb; 
    		10'h2df:	out_reg <= 36'h3eb17cc85; 
    		10'h2e0:	out_reg <= 36'h3ec53ce0f; 
    		10'h2e1:	out_reg <= 36'h3ed87cf9a; 
    		10'h2e2:	out_reg <= 36'h3eeb3d125; 
    		10'h2e3:	out_reg <= 36'h3efd7d2b0; 
    		10'h2e4:	out_reg <= 36'h3f0efd43c; 
    		10'h2e5:	out_reg <= 36'h3f1fbd5c9; 
    		10'h2e6:	out_reg <= 36'h3f2ffd756; 
    		10'h2e7:	out_reg <= 36'h3f3fbd8e3; 
    		10'h2e8:	out_reg <= 36'h3f4ebda70; 
    		10'h2e9:	out_reg <= 36'h3f5d3dbfe; 
    		10'h2ea:	out_reg <= 36'h3f6afdd8d; 
    		10'h2eb:	out_reg <= 36'h3f783df1b; 
    		10'h2ec:	out_reg <= 36'h3f84fe0aa; 
    		10'h2ed:	out_reg <= 36'h3f90fe239; 
    		10'h2ee:	out_reg <= 36'h3f9c3e3c9; 
    		10'h2ef:	out_reg <= 36'h3fa6fe559; 
    		10'h2f0:	out_reg <= 36'h3fb13e6e9; 
    		10'h2f1:	out_reg <= 36'h3fbabe879; 
    		10'h2f2:	out_reg <= 36'h3fc3bea0a; 
    		10'h2f3:	out_reg <= 36'h3fcbfeb9a; 
    		10'h2f4:	out_reg <= 36'h3fd3bed2b; 
    		10'h2f5:	out_reg <= 36'h3fdabeebc; 
    		10'h2f6:	out_reg <= 36'h3fe13f04e; 
    		10'h2f7:	out_reg <= 36'h3fe73f1df; 
    		10'h2f8:	out_reg <= 36'h3fec7f371; 
    		10'h2f9:	out_reg <= 36'h3ff0ff502; 
    		10'h2fa:	out_reg <= 36'h3ff4ff694; 
    		10'h2fb:	out_reg <= 36'h3ff87f826; 
    		10'h2fc:	out_reg <= 36'h3ffb3f9b8; 
    		10'h2fd:	out_reg <= 36'h3ffd3fb4a; 
    		10'h2fe:	out_reg <= 36'h3ffeffcdc; 
    		10'h2ff:	out_reg <= 36'h3fffbfe6e; 
    		10'h300:	out_reg <= 36'h400000000; 
    		10'h301:	out_reg <= 36'h3fff80192; 
    		10'h302:	out_reg <= 36'h3ffec0324; 
    		10'h303:	out_reg <= 36'h3ffd004b6; 
    		10'h304:	out_reg <= 36'h3ffb00648; 
    		10'h305:	out_reg <= 36'h3ff8407da; 
    		10'h306:	out_reg <= 36'h3ff4c096c; 
    		10'h307:	out_reg <= 36'h3ff0c0afe; 
    		10'h308:	out_reg <= 36'h3fec40c8f; 
    		10'h309:	out_reg <= 36'h3fe700e21; 
    		10'h30a:	out_reg <= 36'h3fe100fb2; 
    		10'h30b:	out_reg <= 36'h3fda81144; 
    		10'h30c:	out_reg <= 36'h3fd3812d5; 
    		10'h30d:	out_reg <= 36'h3fcbc1466; 
    		10'h30e:	out_reg <= 36'h3fc3815f6; 
    		10'h30f:	out_reg <= 36'h3fba81787; 
    		10'h310:	out_reg <= 36'h3fb101917; 
    		10'h311:	out_reg <= 36'h3fa6c1aa7; 
    		10'h312:	out_reg <= 36'h3f9c01c37; 
    		10'h313:	out_reg <= 36'h3f90c1dc7; 
    		10'h314:	out_reg <= 36'h3f84c1f56; 
    		10'h315:	out_reg <= 36'h3f78020e5; 
    		10'h316:	out_reg <= 36'h3f6ac2273; 
    		10'h317:	out_reg <= 36'h3f5d02402; 
    		10'h318:	out_reg <= 36'h3f4e82590; 
    		10'h319:	out_reg <= 36'h3f3f8271d; 
    		10'h31a:	out_reg <= 36'h3f2fc28aa; 
    		10'h31b:	out_reg <= 36'h3f1f82a37; 
    		10'h31c:	out_reg <= 36'h3f0ec2bc4; 
    		10'h31d:	out_reg <= 36'h3efd42d50; 
    		10'h31e:	out_reg <= 36'h3eeb02edb; 
    		10'h31f:	out_reg <= 36'h3ed843066; 
    		10'h320:	out_reg <= 36'h3ec5031f1; 
    		10'h321:	out_reg <= 36'h3eb14337b; 
    		10'h322:	out_reg <= 36'h3e9cc3505; 
    		10'h323:	out_reg <= 36'h3e878368e; 
    		10'h324:	out_reg <= 36'h3e71c3817; 
    		10'h325:	out_reg <= 36'h3e5b8399f; 
    		10'h326:	out_reg <= 36'h3e4483b26; 
    		10'h327:	out_reg <= 36'h3e2d03cad; 
    		10'h328:	out_reg <= 36'h3e14c3e33; 
    		10'h329:	out_reg <= 36'h3dfc43fb9; 
    		10'h32a:	out_reg <= 36'h3de2c413e; 
    		10'h32b:	out_reg <= 36'h3dc9042c3; 
    		10'h32c:	out_reg <= 36'h3dae84447; 
    		10'h32d:	out_reg <= 36'h3d93445ca; 
    		10'h32e:	out_reg <= 36'h3d778474d; 
    		10'h32f:	out_reg <= 36'h3d5b448ce; 
    		10'h330:	out_reg <= 36'h3d3e84a50; 
    		10'h331:	out_reg <= 36'h3d2104bd0; 
    		10'h332:	out_reg <= 36'h3d02c4d50; 
    		10'h333:	out_reg <= 36'h3ce444ecf; 
    		10'h334:	out_reg <= 36'h3cc50504d; 
    		10'h335:	out_reg <= 36'h3ca5051ca; 
    		10'h336:	out_reg <= 36'h3c84c5347; 
    		10'h337:	out_reg <= 36'h3c63c54c3; 
    		10'h338:	out_reg <= 36'h3c424563e; 
    		10'h339:	out_reg <= 36'h3c20057b8; 
    		10'h33a:	out_reg <= 36'h3bfd45931; 
    		10'h33b:	out_reg <= 36'h3bda05aaa; 
    		10'h33c:	out_reg <= 36'h3bb605c22; 
    		10'h33d:	out_reg <= 36'h3b9185d98; 
    		10'h33e:	out_reg <= 36'h3b6c85f0e; 
    		10'h33f:	out_reg <= 36'h3b4706083; 
    		10'h340:	out_reg <= 36'h3b20c61f7; 
    		10'h341:	out_reg <= 36'h3afa0636a; 
    		10'h342:	out_reg <= 36'h3ad2c64dc; 
    		10'h343:	out_reg <= 36'h3aaac664d; 
    		10'h344:	out_reg <= 36'h3a82467bd; 
    		10'h345:	out_reg <= 36'h3a594692d; 
    		10'h346:	out_reg <= 36'h3a2fc6a9b; 
    		10'h347:	out_reg <= 36'h3a0586c08; 
    		10'h348:	out_reg <= 36'h39dac6d74; 
    		10'h349:	out_reg <= 36'h39af86edf; 
    		10'h34a:	out_reg <= 36'h3983c7049; 
    		10'h34b:	out_reg <= 36'h3957871b1; 
    		10'h34c:	out_reg <= 36'h392a87319; 
    		10'h34d:	out_reg <= 36'h38fd07480; 
    		10'h34e:	out_reg <= 36'h38cf075e5; 
    		10'h34f:	out_reg <= 36'h38a08774a; 
    		10'h350:	out_reg <= 36'h3871478ad; 
    		10'h351:	out_reg <= 36'h384187a0f; 
    		10'h352:	out_reg <= 36'h381187b70; 
    		10'h353:	out_reg <= 36'h37e0c7cd0; 
    		10'h354:	out_reg <= 36'h37af87e2e; 
    		10'h355:	out_reg <= 36'h377d87f8b; 
    		10'h356:	out_reg <= 36'h374b480e7; 
    		10'h357:	out_reg <= 36'h371848242; 
    		10'h358:	out_reg <= 36'h36e50839c; 
    		10'h359:	out_reg <= 36'h36b1084f4; 
    		10'h35a:	out_reg <= 36'h367c8864b; 
    		10'h35b:	out_reg <= 36'h3647887a1; 
    		10'h35c:	out_reg <= 36'h3612088f5; 
    		10'h35d:	out_reg <= 36'h35dc08a48; 
    		10'h35e:	out_reg <= 36'h35a548b9a; 
    		10'h35f:	out_reg <= 36'h356e48cea; 
    		10'h360:	out_reg <= 36'h3536c8e39; 
    		10'h361:	out_reg <= 36'h34fe88f87; 
    		10'h362:	out_reg <= 36'h34c6090d3; 
    		10'h363:	out_reg <= 36'h348cc921e; 
    		10'h364:	out_reg <= 36'h345349368; 
    		10'h365:	out_reg <= 36'h3419094b0; 
    		10'h366:	out_reg <= 36'h33de895f6; 
    		10'h367:	out_reg <= 36'h33a34973c; 
    		10'h368:	out_reg <= 36'h3367c987f; 
    		10'h369:	out_reg <= 36'h332b899c2; 
    		10'h36a:	out_reg <= 36'h32eec9b02; 
    		10'h36b:	out_reg <= 36'h32b1c9c42; 
    		10'h36c:	out_reg <= 36'h327449d7f; 
    		10'h36d:	out_reg <= 36'h323609ebc; 
    		10'h36e:	out_reg <= 36'h31f789ff6; 
    		10'h36f:	out_reg <= 36'h31b88a12f; 
    		10'h370:	out_reg <= 36'h31790a267; 
    		10'h371:	out_reg <= 36'h3138ca39d; 
    		10'h372:	out_reg <= 36'h30f88a4d2; 
    		10'h373:	out_reg <= 36'h30b78a605; 
    		10'h374:	out_reg <= 36'h30760a736; 
    		10'h375:	out_reg <= 36'h30340a866; 
    		10'h376:	out_reg <= 36'h2ff1ca994; 
    		10'h377:	out_reg <= 36'h2faf0aac0; 
    		10'h378:	out_reg <= 36'h2f6b8abeb; 
    		10'h379:	out_reg <= 36'h2f280ad14; 
    		10'h37a:	out_reg <= 36'h2ee3cae3b; 
    		10'h37b:	out_reg <= 36'h2e9f0af61; 
    		10'h37c:	out_reg <= 36'h2e5a0b085; 
    		10'h37d:	out_reg <= 36'h2e148b1a8; 
    		10'h37e:	out_reg <= 36'h2dce8b2c8; 
    		10'h37f:	out_reg <= 36'h2d880b3e7; 
    		10'h380:	out_reg <= 36'h2d410b504; 
    		10'h381:	out_reg <= 36'h2cf9cb620; 
    		10'h382:	out_reg <= 36'h2cb20b73a; 
    		10'h383:	out_reg <= 36'h2c6a0b852; 
    		10'h384:	out_reg <= 36'h2c214b968; 
    		10'h385:	out_reg <= 36'h2bd84ba7c; 
    		10'h386:	out_reg <= 36'h2b8ecbb8f; 
    		10'h387:	out_reg <= 36'h2b450bca0; 
    		10'h388:	out_reg <= 36'h2afacbdae; 
    		10'h389:	out_reg <= 36'h2ab00bebc; 
    		10'h38a:	out_reg <= 36'h2a650bfc7; 
    		10'h38b:	out_reg <= 36'h2a198c0d0; 
    		10'h38c:	out_reg <= 36'h29cd8c1d8; 
    		10'h38d:	out_reg <= 36'h29814c2de; 
    		10'h38e:	out_reg <= 36'h29348c3e2; 
    		10'h38f:	out_reg <= 36'h28e74c4e3; 
    		10'h390:	out_reg <= 36'h2899cc5e4; 
    		10'h391:	out_reg <= 36'h284bcc6e2; 
    		10'h392:	out_reg <= 36'h27fd8c7de; 
    		10'h393:	out_reg <= 36'h27af0c8d8; 
    		10'h394:	out_reg <= 36'h275fcc9d1; 
    		10'h395:	out_reg <= 36'h27108cac7; 
    		10'h396:	out_reg <= 36'h26c08cbbb; 
    		10'h397:	out_reg <= 36'h26708ccae; 
    		10'h398:	out_reg <= 36'h261fccd9f; 
    		10'h399:	out_reg <= 36'h25cf0ce8d; 
    		10'h39a:	out_reg <= 36'h257d8cf7a; 
    		10'h39b:	out_reg <= 36'h252c0d064; 
    		10'h39c:	out_reg <= 36'h24da0d14d; 
    		10'h39d:	out_reg <= 36'h24878d233; 
    		10'h39e:	out_reg <= 36'h2434cd318; 
    		10'h39f:	out_reg <= 36'h23e1cd3fa; 
    		10'h3a0:	out_reg <= 36'h238e4d4db; 
    		10'h3a1:	out_reg <= 36'h233a8d5b9; 
    		10'h3a2:	out_reg <= 36'h22e68d695; 
    		10'h3a3:	out_reg <= 36'h22920d770; 
    		10'h3a4:	out_reg <= 36'h223d4d848; 
    		10'h3a5:	out_reg <= 36'h21e84d91e; 
    		10'h3a6:	out_reg <= 36'h2192cd9f2; 
    		10'h3a7:	out_reg <= 36'h213d0dac4; 
    		10'h3a8:	out_reg <= 36'h20e70db94; 
    		10'h3a9:	out_reg <= 36'h20908dc61; 
    		10'h3aa:	out_reg <= 36'h2039cdd2d; 
    		10'h3ab:	out_reg <= 36'h1fe2cddf6; 
    		10'h3ac:	out_reg <= 36'h1f8b8debe; 
    		10'h3ad:	out_reg <= 36'h1f340df83; 
    		10'h3ae:	out_reg <= 36'h1edc0e046; 
    		10'h3af:	out_reg <= 36'h1e83ce106; 
    		10'h3b0:	out_reg <= 36'h1e2b4e1c5; 
    		10'h3b1:	out_reg <= 36'h1dd28e282; 
    		10'h3b2:	out_reg <= 36'h1d794e33c; 
    		10'h3b3:	out_reg <= 36'h1d200e3f4; 
    		10'h3b4:	out_reg <= 36'h1cc64e4aa; 
    		10'h3b5:	out_reg <= 36'h1c6c4e55e; 
    		10'h3b6:	out_reg <= 36'h1c124e60f; 
    		10'h3b7:	out_reg <= 36'h1bb7ce6be; 
    		10'h3b8:	out_reg <= 36'h1b5d0e76b; 
    		10'h3b9:	out_reg <= 36'h1b020e816; 
    		10'h3ba:	out_reg <= 36'h1aa6ce8bf; 
    		10'h3bb:	out_reg <= 36'h1a4b4e965; 
    		10'h3bc:	out_reg <= 36'h19ef4ea09; 
    		10'h3bd:	out_reg <= 36'h19934eaab; 
    		10'h3be:	out_reg <= 36'h19370eb4b; 
    		10'h3bf:	out_reg <= 36'h18da8ebe8; 
    		10'h3c0:	out_reg <= 36'h187dcec83; 
    		10'h3c1:	out_reg <= 36'h1820ced1c; 
    		10'h3c2:	out_reg <= 36'h17c38edb2; 
    		10'h3c3:	out_reg <= 36'h17660ee46; 
    		10'h3c4:	out_reg <= 36'h17088eed8; 
    		10'h3c5:	out_reg <= 36'h16aa8ef68; 
    		10'h3c6:	out_reg <= 36'h164c4eff5; 
    		10'h3c7:	out_reg <= 36'h15ee0f080; 
    		10'h3c8:	out_reg <= 36'h158f8f109; 
    		10'h3c9:	out_reg <= 36'h1530cf18f; 
    		10'h3ca:	out_reg <= 36'h14d1cf213; 
    		10'h3cb:	out_reg <= 36'h14728f294; 
    		10'h3cc:	out_reg <= 36'h14134f314; 
    		10'h3cd:	out_reg <= 36'h13b3cf391; 
    		10'h3ce:	out_reg <= 36'h13540f40b; 
    		10'h3cf:	out_reg <= 36'h12f40f484; 
    		10'h3d0:	out_reg <= 36'h12940f4fa; 
    		10'h3d1:	out_reg <= 36'h12338f56d; 
    		10'h3d2:	out_reg <= 36'h11d34f5de; 
    		10'h3d3:	out_reg <= 36'h11728f64d; 
    		10'h3d4:	out_reg <= 36'h1111cf6ba; 
    		10'h3d5:	out_reg <= 36'h10b0cf724; 
    		10'h3d6:	out_reg <= 36'h104f8f78b; 
    		10'h3d7:	out_reg <= 36'h0fee4f7f1; 
    		10'h3d8:	out_reg <= 36'h0f8ccf853; 
    		10'h3d9:	out_reg <= 36'h0f2b4f8b4; 
    		10'h3da:	out_reg <= 36'h0ec98f912; 
    		10'h3db:	out_reg <= 36'h0e67cf96e; 
    		10'h3dc:	out_reg <= 36'h0e05cf9c7; 
    		10'h3dd:	out_reg <= 36'h0da38fa1e; 
    		10'h3de:	out_reg <= 36'h0d414fa73; 
    		10'h3df:	out_reg <= 36'h0cdecfac5; 
    		10'h3e0:	out_reg <= 36'h0c7c4fb14; 
    		10'h3e1:	out_reg <= 36'h0c198fb61; 
    		10'h3e2:	out_reg <= 36'h0bb6cfbac; 
    		10'h3e3:	out_reg <= 36'h0b540fbf5; 
    		10'h3e4:	out_reg <= 36'h0af10fc3b; 
    		10'h3e5:	out_reg <= 36'h0a8dcfc7e; 
    		10'h3e6:	out_reg <= 36'h0a2a8fcbf; 
    		10'h3e7:	out_reg <= 36'h09c74fcfe; 
    		10'h3e8:	out_reg <= 36'h09640fd3a; 
    		10'h3e9:	out_reg <= 36'h09008fd74; 
    		10'h3ea:	out_reg <= 36'h089ccfdab; 
    		10'h3eb:	out_reg <= 36'h08394fde0; 
    		10'h3ec:	out_reg <= 36'h07d58fe13; 
    		10'h3ed:	out_reg <= 36'h0771cfe43; 
    		10'h3ee:	out_reg <= 36'h070dcfe70; 
    		10'h3ef:	out_reg <= 36'h06a9cfe9b; 
    		10'h3f0:	out_reg <= 36'h0645cfec4; 
    		10'h3f1:	out_reg <= 36'h05e1cfeea; 
    		10'h3f2:	out_reg <= 36'h057d8ff0e; 
    		10'h3f3:	out_reg <= 36'h05198ff2f; 
    		10'h3f4:	out_reg <= 36'h04b54ff4e; 
    		10'h3f5:	out_reg <= 36'h04510ff6a; 
    		10'h3f6:	out_reg <= 36'h03ec8ff84; 
    		10'h3f7:	out_reg <= 36'h03884ff9c; 
    		10'h3f8:	out_reg <= 36'h0323cffb1; 
    		10'h3f9:	out_reg <= 36'h02bf8ffc3; 
    		10'h3fa:	out_reg <= 36'h025b0ffd3; 
    		10'h3fb:	out_reg <= 36'h01f68ffe1; 
    		10'h3fc:	out_reg <= 36'h01920ffec; 
    		10'h3fd:	out_reg <= 36'h012d8fff4; 
    		10'h3fe:	out_reg <= 36'h00c90fffb; 
    		10'h3ff:	out_reg <= 36'h00648fffe; 
    		default: out_reg <= 0;
    	endcase
    end
end
endgenerate

endmodule

